`timescale 1ns / 1ps
`default_nettype none
//
// RISu64
// Copyright 2022 Wenting Zhang
//
// Permission is hereby granted, free of charge, to any person obtaining a copy
// of this software and associated documentation files (the "Software"), to deal
// in the Software without restriction, including without limitation the rights
// to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
// copies of the Software, and to permit persons to whom the Software is
// furnished to do so, subject to the following conditions:
//
// The above copyright notice and this permission notice shall be included in
// all copies or substantial portions of the Software.
//
// THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
// IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
// FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
// AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
// LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
// OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
// SOFTWARE.
//
`include "defines.vh"

module ix(
    input  wire         clk,
    input  wire         rst,
    input  wire         pipe_flush,
    // Register file interface
    output wire [4:0]   rf_rsrc0,
    input  wire [63:0]  rf_rdata0,
    output wire [4:0]   rf_rsrc1,
    input  wire [63:0]  rf_rdata1,
    output wire [4:0]   rf_rsrc2,
    input  wire [63:0]  rf_rdata2,
    output wire [4:0]   rf_rsrc3,
    input  wire [63:0]  rf_rdata3,
    // IX interface
    input  wire [247:0] dec0_ix_bundle,
    input  wire         dec0_ix_valid,
    output wire         dec0_ix_ready,
    input  wire [247:0] dec1_ix_bundle,
    input  wire         dec1_ix_valid,
    output wire         dec1_ix_ready,
    // FU interfaces
    // To integer pipe 0
    output reg  [63:0]  ix_ip0_pc,
    output reg  [4:0]   ix_ip0_dst,
    output reg          ix_ip0_wb_en,
    output reg  [3:0]   ix_ip0_op,
    output reg          ix_ip0_option,
    output reg          ix_ip0_truncate,
    output reg  [1:0]   ix_ip0_br_type,
    output reg          ix_ip0_br_neg,
    output reg  [63:0]  ix_ip0_br_base,
    output reg  [20:0]  ix_ip0_br_offset,
    output reg          ix_ip0_br_is_call,
    output reg          ix_ip0_br_is_ret,
    output reg  [63:0]  ix_ip0_operand1,
    output reg  [63:0]  ix_ip0_operand2,
    output reg          ix_ip0_bp,
    output reg  [1:0]   ix_ip0_bp_track,
    output reg  [63:0]  ix_ip0_bt,
    output reg          ix_ip0_valid,
    input  wire         ix_ip0_ready,
    // Hazard detection & Bypassing
    input  wire [63:0]  ip0_ix_forwarding,
    input  wire [4:0]   ip0_wb_dst,
    input  wire [63:0]  ip0_wb_result,
    input  wire         ip0_wb_wb_en,
    input  wire         ip0_wb_valid,
    // To integer pipe 1
    output reg  [63:0]  ix_ip1_pc,
    output reg  [4:0]   ix_ip1_dst,
    output reg          ix_ip1_wb_en,
    output reg  [3:0]   ix_ip1_op,
    output reg          ix_ip1_option,
    output reg          ix_ip1_truncate,
    output reg  [1:0]   ix_ip1_br_type,
    output reg          ix_ip1_br_neg,
    output reg  [63:0]  ix_ip1_br_base,
    output reg  [20:0]  ix_ip1_br_offset,
    output reg          ix_ip1_br_is_call,
    output reg          ix_ip1_br_is_ret,
    output reg  [63:0]  ix_ip1_operand1,
    output reg  [63:0]  ix_ip1_operand2,
    output reg          ix_ip1_bp,
    output reg  [1:0]   ix_ip1_bp_track,
    output reg  [63:0]  ix_ip1_bt,
    output reg          ix_ip1_speculate,
    output reg          ix_ip1_valid,
    input  wire         ix_ip1_ready,
    // Hazard detection & Bypassing
    input  wire [63:0]  ip1_ix_forwarding,
    input  wire [4:0]   ip1_wb_dst,
    input  wire [63:0]  ip1_wb_result,
    input  wire         ip1_wb_wb_en,
    input  wire         ip1_wb_valid,
    // To load/ store pipe
    output reg  [63:0]  ix_lsp_pc,
    output reg  [4:0]   ix_lsp_dst,
    output reg          ix_lsp_wb_en,
    output reg  [63:0]  ix_lsp_base,
    output reg  [11:0]  ix_lsp_offset,
    output reg  [63:0]  ix_lsp_source,
    output reg          ix_lsp_mem_sign,
    output reg  [1:0]   ix_lsp_mem_width,
    output reg          ix_lsp_speculate,
    output reg          ix_lsp_valid,
    input  wire         ix_lsp_ready,
    input  wire         lsp_unaligned_load,
    input  wire         lsp_unaligned_store,
    input  wire [63:0]  lsp_unaligned_epc,
    // Hazard detection & Bypassing
    input  wire         lsp_ix_mem_busy,
    input  wire         lsp_ix_mem_wb_en,
    input  wire [4:0]   lsp_ix_mem_dst,
    input  wire [63:0]  lsp_ix_mem_result,
    input  wire         lsp_ix_mem_result_valid,
    input  wire [4:0]   lsp_wb_dst,
    input  wire [63:0]  lsp_wb_result,
    input  wire         lsp_wb_wb_en,
    input  wire         lsp_wb_valid,
    // To muldiv unit
    output reg  [63:0]  ix_md_pc,
    output reg  [4:0]   ix_md_dst,
    output reg  [63:0]  ix_md_operand1,
    output reg  [63:0]  ix_md_operand2,
    output reg  [2:0]   ix_md_md_op,
    output reg          ix_md_muldiv,
    output reg          ix_md_speculate,
    output reg          ix_md_valid,
    input  wire         ix_md_ready,
    // Hazard detection
    input  wire [4:0]   md_ix_dst,
    input  wire         md_ix_active,
    // To trap unit
    output reg  [63:0]  ix_trap_pc,
    output reg  [4:0]   ix_trap_dst,
    output reg  [1:0]   ix_trap_csr_op,
    output reg  [11:0]  ix_trap_csr_id,
    output reg  [63:0]  ix_trap_csr_opr,
    output reg          ix_trap_mret,
    output reg          ix_trap_int,
    output reg          ix_trap_intexc,
    output reg  [3:0]   ix_trap_cause,
    output reg          ix_trap_valid,
    input  wire         ix_trap_ready,
    input  wire [15:0]  trap_ix_ip,
    // From WB
    input  wire [63:0]  wb_ix_buf_value,
    input  wire [4:0]   wb_ix_buf_dst,
    input  wire         wb_ix_buf_valid,
    // MMU
    input  wire         mmu_load_page_fault,
    input  wire         mmu_store_page_fault,
    input  wire [63:0]  mmu_fault_epc,
    output wire         ix_mmu_tlb_flush_req,
    // Fence I
    output reg          im_invalidate_req,
    input  wire         im_invalidate_resp,
    output reg          dm_flush_req,
    input  wire         dm_flush_resp,
    output reg          ix_if_pc_override,
    output reg  [63:0]  ix_if_new_pc
);

    // Unbundle signals
    wire [63:0] dec0_ix_pc;
    wire        dec0_ix_bp;
    wire [1:0]  dec0_ix_bp_track;
    wire [63:0] dec0_ix_bt;
    wire [3:0]  dec0_ix_op;
    wire        dec0_ix_option;
    wire        dec0_ix_truncate;
    wire [1:0]  dec0_ix_br_type;
    wire        dec0_ix_br_neg;
    wire        dec0_ix_br_base_src;
    wire        dec0_ix_br_inj_pc;
    wire        dec0_ix_br_is_call;
    wire        dec0_ix_br_is_ret;
    wire        dec0_ix_mem_sign;
    wire [1:0]  dec0_ix_mem_width;
    wire [1:0]  dec0_ix_csr_op;
    wire        dec0_ix_mret;
    wire        dec0_ix_intr;
    wire [3:0]  dec0_ix_cause;
    wire [2:0]  dec0_ix_md_op;
    wire        dec0_ix_muldiv;
    wire [2:0]  dec0_ix_op_type;
    wire [1:0]  dec0_ix_operand1;
    wire [1:0]  dec0_ix_operand2;
    wire [63:0] dec0_ix_imm;
    wire        dec0_ix_legal;
    wire        dec0_ix_wb_en;
    wire [4:0]  dec0_ix_rs1;
    wire [4:0]  dec0_ix_rs2;
    wire [4:0]  dec0_ix_rd;
    wire        dec0_ix_fencei;

    wire [63:0] dec1_ix_pc;
    wire        dec1_ix_bp;
    wire [1:0]  dec1_ix_bp_track;
    wire [63:0] dec1_ix_bt;
    wire [3:0]  dec1_ix_op;
    wire        dec1_ix_option;
    wire        dec1_ix_truncate;
    wire [1:0]  dec1_ix_br_type;
    wire        dec1_ix_br_neg;
    wire        dec1_ix_br_base_src;
    wire        dec1_ix_br_inj_pc;
    wire        dec1_ix_br_is_call;
    wire        dec1_ix_br_is_ret;
    wire        dec1_ix_mem_sign;
    wire [1:0]  dec1_ix_mem_width;
    wire [1:0]  dec1_ix_csr_op;
    wire        dec1_ix_mret;
    wire        dec1_ix_intr;
    wire [3:0]  dec1_ix_cause;
    wire [2:0]  dec1_ix_md_op;
    wire        dec1_ix_muldiv;
    wire [2:0]  dec1_ix_op_type;
    wire [1:0]  dec1_ix_operand1;
    wire [1:0]  dec1_ix_operand2;
    wire [63:0] dec1_ix_imm;
    wire        dec1_ix_legal;
    wire        dec1_ix_wb_en;
    wire [4:0]  dec1_ix_rs1;
    wire [4:0]  dec1_ix_rs2;
    wire [4:0]  dec1_ix_rd;
    wire        dec1_ix_fencei;

    assign {
        dec0_ix_pc,
        dec0_ix_bp,
        dec0_ix_bp_track,
        dec0_ix_bt,
        dec0_ix_op,
        dec0_ix_option,
        dec0_ix_truncate,
        dec0_ix_br_type,
        dec0_ix_br_neg,
        dec0_ix_br_base_src,
        dec0_ix_br_inj_pc,
        dec0_ix_br_is_call,
        dec0_ix_br_is_ret,
        dec0_ix_mem_sign,
        dec0_ix_mem_width,
        dec0_ix_csr_op,
        dec0_ix_mret,
        dec0_ix_intr,
        dec0_ix_cause,
        dec0_ix_md_op,
        dec0_ix_muldiv,
        dec0_ix_op_type,
        dec0_ix_operand1,
        dec0_ix_operand2,
        dec0_ix_imm,
        dec0_ix_legal,
        dec0_ix_wb_en,
        dec0_ix_rs1,
        dec0_ix_rs2,
        dec0_ix_rd,
        dec0_ix_fencei} = dec0_ix_bundle;
    
    assign {
        dec1_ix_pc,
        dec1_ix_bp,
        dec1_ix_bp_track,
        dec1_ix_bt,
        dec1_ix_op,
        dec1_ix_option,
        dec1_ix_truncate,
        dec1_ix_br_type,
        dec1_ix_br_neg,
        dec1_ix_br_base_src,
        dec1_ix_br_inj_pc,
        dec1_ix_br_is_call,
        dec1_ix_br_is_ret,
        dec1_ix_mem_sign,
        dec1_ix_mem_width,
        dec1_ix_csr_op,
        dec1_ix_mret,
        dec1_ix_intr,
        dec1_ix_cause,
        dec1_ix_md_op,
        dec1_ix_muldiv,
        dec1_ix_op_type,
        dec1_ix_operand1,
        dec1_ix_operand2,
        dec1_ix_imm,
        dec1_ix_legal,
        dec1_ix_wb_en,
        dec1_ix_rs1,
        dec1_ix_rs2,
        dec1_ix_rd,
        dec1_ix_fencei} = dec1_ix_bundle;

    // Hazard detection
    assign rf_rsrc0 = dec0_ix_rs1;
    assign rf_rsrc1 = dec0_ix_rs2;
    assign rf_rsrc2 = dec1_ix_rs1;
    assign rf_rsrc3 = dec1_ix_rs2;
    wire [4:0] rf_rsrc [0:3];
    assign rf_rsrc[0] = rf_rsrc0;
    assign rf_rsrc[1] = rf_rsrc1;
    assign rf_rsrc[2] = rf_rsrc2;
    assign rf_rsrc[3] = rf_rsrc3;
    wire [63:0] rf_rdata [0:3];
    assign rf_rdata[0] = rf_rdata0;
    assign rf_rdata[1] = rf_rdata1;
    assign rf_rdata[2] = rf_rdata2;
    assign rf_rdata[3] = rf_rdata3;
    reg [0:0] rs_ready [0:3];
    reg [63:0] rs_val [0:3];
    wire ip0_ex_ixstalled = ix_ip0_valid && !ix_ip0_ready && ix_ip0_wb_en;
    wire ip0_ex_active = ix_ip0_valid && ix_ip0_ready && ix_ip0_wb_en;
    wire ip0_wb_active = ip0_wb_valid && ip0_wb_wb_en;
    wire ip1_ex_ixstalled = ix_ip1_valid && !ix_ip1_ready && ix_ip1_wb_en;
    wire ip1_ex_active = ix_ip1_valid && ix_ip1_ready && ix_ip1_wb_en;
    wire ip1_wb_active = ip1_wb_valid && ip1_wb_wb_en;
    wire lsp_ag_active = ix_lsp_valid;
    wire lsp_mem_active = lsp_ix_mem_busy;
    wire lsp_wb_active = lsp_wb_valid && lsp_wb_wb_en;
    /* verilator lint_off UNUSED */
    reg dbg_stl_ip0 [0:3];
    reg dbg_stl_ip1 [0:3];
    reg dbg_stl_lag [0:3];
    reg dbg_stl_lma [0:3];
    reg dbg_stl_mdi [0:3];
    reg dbg_stl_mda [0:3];
    /* verilator lint_on UNUSED */
    genvar i;
    generate
        for (i = 0; i < 4; i = i + 1) begin
            always @(*) begin
                dbg_stl_ip0[i] = 1'b0;
                dbg_stl_ip1[i] = 1'b0;
                dbg_stl_lag[i] = 1'b0;
                dbg_stl_lma[i] = 1'b0;
                dbg_stl_mdi[i] = 1'b0;
                dbg_stl_mda[i] = 1'b0;

                rs_ready[i] = 1'b1;
                // Register read
                rs_val[i] = (rf_rsrc[i] == 5'd0) ? (64'd0) : rf_rdata[i];

                // Must be from late to early in case there are WAW dependencies
                // The ordering only applies to within the FU: inter-FU
                // (non-deterministic) WAW is handled previously.

                // Forwarding point: WB buffer
                if (wb_ix_buf_valid && (wb_ix_buf_dst == rf_rsrc[i])) begin
                    rs_ready[i] = 1'b1;
                    rs_val[i] = wb_ix_buf_value;
                end
                // Forwarding point: IP0 writeback
                if (ip0_wb_active && (ip0_wb_dst == rf_rsrc[i])) begin
                    rs_ready[i] = 1'b1;
                    rs_val[i] = ip0_wb_result;
                end
                if (ip1_wb_active && (ip1_wb_dst == rf_rsrc[i])) begin
                    rs_ready[i] = 1'b1;
                    rs_val[i] = ip1_wb_result;
                end
                // Forwarding point: IP1 execution
                if (ip0_ex_active && (ix_ip0_dst == rf_rsrc[i])) begin
                    rs_ready[i] = 1'b1;
                    rs_val[i] = ip0_ix_forwarding;
                end
                if (ip1_ex_active && (ix_ip1_dst == rf_rsrc[i])) begin
                    rs_ready[i] = 1'b1;
                    rs_val[i] = ip1_ix_forwarding;
                end
                // Stall point: IP execution not accepted
                if (ip0_ex_ixstalled && (ix_ip0_dst == rf_rsrc[i])) begin
                    rs_ready[i] = 1'b0;
                    dbg_stl_ip0[i] = 1'b1;
                end
                if (ip1_ex_ixstalled && (ix_ip1_dst == rf_rsrc[i])) begin
                    rs_ready[i] = 1'b0;
                    dbg_stl_ip1[i] = 1'b1;
                end

                // Forwarding point: LSP writeback
                if (lsp_wb_active && (lsp_wb_dst == rf_rsrc[i])) begin
                    rs_ready[i] = 1'b1;
                    rs_val[i] = lsp_wb_result;
                end
                // Stall point: LSP memory access active
                if (lsp_ix_mem_wb_en && (lsp_ix_mem_dst == rf_rsrc[i])) begin
                    rs_ready[i] = 1'b0;
                    dbg_stl_lma[i] = 1'b1;
                end
                // Forwarding point: LSP readout
                `ifdef ENABLE_MEM_FORWARING
                if (lsp_ix_mem_wb_en && (lsp_ix_mem_dst == rf_rsrc[i]) &&
                        lsp_ix_mem_result_valid) begin
                    rs_ready[i] = 1'b1;
                    rs_val[i] = lsp_ix_mem_result;
                end
                `endif
                // Stall point: LSP address generation
                if (lsp_ag_active && ix_lsp_wb_en &&
                        (ix_lsp_dst == rf_rsrc[i])) begin
                    rs_ready[i] = 1'b0;
                    dbg_stl_lag[i] = 1'b1;
                end
                // Stall point: MD issue
                if (ix_md_valid && (ix_md_dst == rf_rsrc[i])) begin
                    rs_ready[i] = 1'b0;
                    dbg_stl_mdi[i] = 1'b1;
                end
                // Stall point: MD active
                if (md_ix_active && (md_ix_dst == rf_rsrc[i])) begin
                    rs_ready[i] = 1'b0;
                    dbg_stl_mda[i] = 1'b1;
                end

                // Always override to 0 in case write to 0 forwarding is valid
                if (rf_rsrc[i] == 5'd0) begin
                    rs_ready[i] = 1'b1;
                    rs_val[i] = 64'd0;
                end
            end
        end
    endgenerate

    // WAW hazard
    // TODO: If WB is accepted this cycle OR will be accepted next cycle,
    // then it's not a hazard
    wire waw_from_ip0_dec0 = (!dec0_ix_wb_en) ||
            ((!ip0_wb_active || (ip0_wb_dst != dec0_ix_rd)) &&
            (!ip0_ex_active || (ix_ip0_dst != dec0_ix_rd)) &&
            (!ip0_ex_ixstalled || (ix_ip0_dst != dec0_ix_rd)));
    wire waw_from_ip0_dec1 = (!dec1_ix_wb_en) ||
            ((!ip0_wb_active || (ip0_wb_dst != dec1_ix_rd)) &&
            (!ip0_ex_active || (ix_ip0_dst != dec1_ix_rd)) &&
            (!ip0_ex_ixstalled || (ix_ip0_dst != dec1_ix_rd)));
    wire waw_from_ip1_dec0 = (!dec0_ix_wb_en) ||
            ((!ip1_wb_active || (ip1_wb_dst != dec0_ix_rd)) &&
            (!ip1_ex_active || (ix_ip1_dst != dec0_ix_rd)) &&
            (!ip1_ex_ixstalled || (ix_ip1_dst != dec0_ix_rd)));
    wire waw_from_ip1_dec1 = (!dec1_ix_wb_en) ||
            ((!ip1_wb_active || (ip1_wb_dst != dec1_ix_rd)) &&
            (!ip1_ex_active || (ix_ip1_dst != dec1_ix_rd)) &&
            (!ip1_ex_ixstalled || (ix_ip1_dst != dec1_ix_rd)));
    wire waw_from_ip_dec0 = waw_from_ip0_dec0 && waw_from_ip1_dec0;
    wire waw_from_ip_dec1 = waw_from_ip0_dec1 && waw_from_ip1_dec1;
    // Warning: this doesn't check the case where LSP is ready for WB.
    // This is creates an edge case where is a load instruction destination is
    // also used for jal target register, and MD happens to be active for two
    // cycles (doesn't currently possible), a WAW condition happens.
    // When this ever becomes possible, WB stage needs provision to fix this.
    wire waw_from_lsp_dec0 =
            (!lsp_ix_mem_wb_en || (lsp_ix_mem_dst != dec0_ix_rd)) &&
            (!lsp_ag_active || !ix_lsp_wb_en || (ix_lsp_dst != dec0_ix_rd));
    wire waw_from_lsp_dec1 =
            (!lsp_ix_mem_wb_en || (lsp_ix_mem_dst != dec1_ix_rd)) &&
            (!lsp_ag_active || !ix_lsp_wb_en || (ix_lsp_dst != dec1_ix_rd));
    wire waw_from_md_dec0 = (!ix_md_valid || (ix_md_dst != dec0_ix_rd)) &&
            (!md_ix_active || (md_ix_dst != dec0_ix_rd));
    wire waw_from_md_dec1 = (!ix_md_valid || (ix_md_dst != dec1_ix_rd)) &&
            (!md_ix_active || (md_ix_dst != dec1_ix_rd));
    // For LSP: It's only going to be faster than MD, only check md
    wire waw_lsp_dec0 = waw_from_ip_dec0 && waw_from_md_dec0;
    wire waw_lsp_dec1 = waw_from_ip_dec1 && waw_from_md_dec1;
    // For IP: It need to protect against LSP and MD
    wire waw_ip_dec0 = waw_from_lsp_dec0 && waw_from_md_dec0;
    wire waw_ip_dec1 = waw_from_lsp_dec1 && waw_from_md_dec1;
    // For MD: It need to protect against only LSP
    wire waw_md_dec0 = waw_from_lsp_dec0;
    wire waw_md_dec1 = waw_from_lsp_dec1;

    wire operand1_dec0_ready = (dec0_ix_operand1 == `D_OPR1_RS1) ? rs_ready[0] : 1'b1;
    wire operand2_dec0_ready = (dec0_ix_operand2 == `D_OPR2_RS2) ? rs_ready[1] : 1'b1;
    wire operand1_dec1_ready = (dec1_ix_operand1 == `D_OPR1_RS1) ? rs_ready[2] : 1'b1;
    wire operand2_dec1_ready = (dec1_ix_operand2 == `D_OPR2_RS2) ? rs_ready[3] : 1'b1;

    wire [63:0] operand1_dec0_value = ((dec0_ix_operand1 == `D_OPR1_PC) ||
            (dec0_ix_br_inj_pc)) ? (dec0_ix_pc) :
            (dec0_ix_operand1 == `D_OPR1_RS1) ? (rs_val[0]) :
            (dec0_ix_operand1 == `D_OPR1_ZERO) ? (64'd0) :
            (dec0_ix_operand1 == `D_OPR1_ZIMM) ? ({59'd0, dec0_ix_rs1}) : (64'bx);
    wire [63:0] operand2_dec0_value =
            (dec0_ix_operand2 == `D_OPR2_RS2) ? (rs_val[1]) :
            (dec0_ix_operand2 == `D_OPR2_IMM) ? (dec0_ix_imm) :
            (dec0_ix_operand2 == `D_OPR2_4) ? (64'd4) : (64'bx);
    wire [63:0] operand1_dec1_value = ((dec1_ix_operand1 == `D_OPR1_PC) ||
            (dec1_ix_br_inj_pc)) ? (dec1_ix_pc) :
            (dec1_ix_operand1 == `D_OPR1_RS1) ? (rs_val[2]) :
            (dec1_ix_operand1 == `D_OPR1_ZERO) ? (64'd0) :
            (dec1_ix_operand1 == `D_OPR1_ZIMM) ? ({59'd0, dec1_ix_rs1}) : (64'bx);
    wire [63:0] operand2_dec1_value =
            (dec1_ix_operand2 == `D_OPR2_RS2) ? (rs_val[3]) :
            (dec1_ix_operand2 == `D_OPR2_IMM) ? (dec1_ix_imm) :
            (dec1_ix_operand2 == `D_OPR2_4) ? (64'd4) : (64'bx);

    wire [63:0] br_base_dec0 = (dec0_ix_br_base_src == `BB_PC) ? (dec0_ix_pc) :
            (rs_val[0]);
    wire [63:0] br_base_dec1 = (dec1_ix_br_base_src == `BB_PC) ? (dec1_ix_pc) :
            (rs_val[2]);

    // Trap instruction also blocks all proceeding instructions
    reg trap_ongoing;
    wire int_pending = (trap_ix_ip != 16'd0);
    wire lsp_fault = lsp_unaligned_load || lsp_unaligned_store;
    wire mmu_fault = mmu_load_page_fault || mmu_store_page_fault;
    wire exc_pending = lsp_fault || mmu_fault;
    wire ix_dec0_opr_ready = operand1_dec0_ready && operand2_dec0_ready;
    wire ix_dec1_opr_ready = operand1_dec1_ready && operand2_dec1_ready;
    wire lsp_req_pending = ix_lsp_valid;
    wire md_req_pending = ix_md_valid;
    wire ix_issue_common = !pipe_flush && !trap_ongoing && !int_pending &&
            !exc_pending;
    wire dec0_is_int = (dec0_ix_op_type == `OT_INT);
    wire dec1_is_int = (dec1_ix_op_type == `OT_INT);
    wire dec0_is_ls = ((dec0_ix_op_type == `OT_LOAD) || (dec0_ix_op_type == `OT_STORE));
    wire dec1_is_ls = ((dec1_ix_op_type == `OT_LOAD) || (dec1_ix_op_type == `OT_STORE));
    wire dec1_is_load = (dec1_ix_op_type == `OT_LOAD);
    wire dec0_is_md = (dec0_ix_op_type == `OT_MULDIV);
    wire dec1_is_md = (dec1_ix_op_type == `OT_MULDIV);
    wire dec0_is_branch = (dec0_ix_op_type == `OT_BRANCH);
    wire dec1_is_branch = (dec1_ix_op_type == `OT_BRANCH);
    wire dec0_is_trap = (dec0_ix_op_type == `OT_TRAP);
    wire dec0_is_fence = (dec0_ix_op_type == `OT_FENCE);

    // Inter-dependency check:
    // 1. Both decoded instructions are valid
    // 2. They should not write to the same register
    // 3. INST0 should not write to one of the source of INST1
    wire ix_interdep_check = dec0_ix_valid && dec1_ix_valid &&
            ((dec0_ix_rd != dec1_ix_rd) || !(dec0_ix_wb_en && dec1_ix_wb_en)) &&
            (!dec0_ix_wb_en || (
                ((dec0_ix_rd != dec1_ix_rs1) || (dec1_ix_operand1 != `D_OPR1_RS1)) &&
                ((dec0_ix_rd != dec1_ix_rs2) || (dec1_ix_operand2 != `D_OPR2_RS2)))) &&
            (!dec0_is_branch || dec1_is_int || dec1_is_md || dec1_is_load);
    // Issue logic

    wire ix_fenced_done = !(lsp_ag_active || lsp_mem_active || lsp_wb_active);
    reg ix_fencei_done = 1'b0;
    // Wait for integer pipe to finish
    wire ix_ibarrier_done = !(ip0_ex_ixstalled || ip0_ex_active || ip0_wb_active);
    // Barrier for waiting for in-flight instructions to complete
    wire ix_barrier_done = ix_fenced_done && ix_ibarrier_done;

    reg ix_issue_ip0_dec0;
    reg ix_issue_ip1_dec1;
    reg ix_issue_lsp_dec0;
    reg ix_issue_lsp_dec1;
    reg ix_issue_md_dec0;
    reg ix_issue_md_dec1;
    reg ix_issue_trap;
    reg ix_fence_done;

    reg ix_issue_dec0;
    reg ix_issue_dec1;
    always @(*) begin
        ix_issue_ip0_dec0 = 0;
        ix_issue_ip1_dec1 = 0;
        ix_issue_lsp_dec0 = 0;
        ix_issue_lsp_dec1 = 0;
        ix_issue_md_dec0 = 0;
        ix_issue_md_dec1 = 0;
        ix_issue_trap = 0;
        ix_fence_done = 0;
        ix_issue_dec0 = 0;
        ix_issue_dec1 = 0;
        if (ix_issue_common && dec0_ix_valid && ix_dec0_opr_ready) begin
            // Trap and fence are not handled here
            if (dec0_is_int && waw_ip_dec0 && ix_ip0_ready) begin
                ix_issue_dec0 = 1;
                ix_issue_ip0_dec0 = 1;
            end
            if (dec0_is_branch && waw_ip_dec0 && ix_ip0_ready &&
                    !lsp_req_pending && !md_req_pending) begin
                ix_issue_dec0 = 1;
                ix_issue_ip0_dec0 = 1;
            end
            else if (dec0_is_ls && waw_lsp_dec0 && ix_lsp_ready) begin
                ix_issue_dec0 = 1;
                ix_issue_lsp_dec0 = 1;
            end
            else if (dec0_is_md && waw_md_dec0 && ix_md_ready) begin
                ix_issue_dec0 = 1;
                ix_issue_md_dec0 = 1;
            end
            else if (dec0_is_trap && !trap_ongoing && ix_barrier_done) begin
                ix_issue_dec0 = 1;
                ix_issue_trap = 1;
            end
            else if (dec0_is_fence && ix_fenced_done &&
                    (!dec0_ix_fencei || ix_fencei_done)) begin
                ix_issue_dec0 = 1;
                ix_fence_done = 1;
            end

            if (ix_issue_dec0 && ix_interdep_check && ix_dec1_opr_ready) begin
                // Can issue the second one?
                if (dec1_is_int && waw_ip_dec1 && ix_ip1_ready) begin
                    ix_issue_dec1 = 1;
                    ix_issue_ip1_dec1 = 1;
                end
                else if (dec1_is_branch && waw_ip_dec1 && ix_ip1_ready &&
                        !lsp_req_pending && !md_req_pending) begin
                    ix_issue_dec1 = 1;
                    ix_issue_ip1_dec1 = 1;
                end
                else if (dec1_is_ls && waw_lsp_dec1 && !dec0_is_ls && ix_lsp_ready) begin
                    ix_issue_dec1 = 1;
                    ix_issue_lsp_dec1 = 1;
                end
                else if (dec1_is_md && waw_md_dec1 && !dec0_is_md && ix_md_ready) begin
                    ix_issue_dec1 = 1;
                    ix_issue_md_dec1 = 1;
                end
            end
        end
    end

    // TODO: Implement actual sfence.vma support
    assign ix_mmu_tlb_flush_req = ix_fence_done;

    wire ix_issue_ip0 = ix_issue_ip0_dec0;
    wire ix_issue_ip1 = ix_issue_ip1_dec1;
    wire ix_issue_lsp = ix_issue_lsp_dec0 || ix_issue_lsp_dec1;
    wire ix_issue_md = ix_issue_md_dec0 || ix_issue_md_dec1;

    wire ix_stall = dec0_ix_valid && !ix_issue_dec0 && !pipe_flush;
    assign dec0_ix_ready = !rst && !ix_stall;
    assign dec1_ix_ready = !rst && !ix_stall && ix_issue_dec1;

    reg [63:0] dbg_cntr_fe_stall;
    reg [63:0] dbg_cntr_no_issue;
    reg [63:0] dbg_cntr_one_issue;
    reg [63:0] dbg_cntr_dep_fail;
    reg [63:0] dbg_cntr_dep_raw;
    reg [63:0] dbg_cntr_dep_waw;
    reg [63:0] dbg_cntr_str_brbr;
    reg [63:0] dbg_cntr_str_brls;
    reg [63:0] dbg_cntr_str_brother;
    reg [63:0] dbg_cntr_dual_issue;
    always @(posedge clk) begin
        if (ix_issue_dec0 ^ ix_issue_dec1)
            dbg_cntr_one_issue <= dbg_cntr_one_issue + 1;
        else if (ix_issue_dec0 && ix_issue_dec1)
            dbg_cntr_dual_issue <= dbg_cntr_dual_issue + 1;
        else
            dbg_cntr_no_issue <= dbg_cntr_no_issue + 1;
        if (!dec0_ix_valid)
            dbg_cntr_fe_stall <= dbg_cntr_fe_stall + 1;
        if (dbg_cntr_one_issue && dec1_ix_valid && !ix_interdep_check) begin
            dbg_cntr_dep_fail <= dbg_cntr_dep_fail + 1;
            if (dec0_ix_wb_en && (
            ((dec0_ix_rd == dec1_ix_rs1) && (dec1_ix_operand1 == `D_OPR1_RS1)) ||
            ((dec0_ix_rd == dec1_ix_rs2) && (dec1_ix_operand2 == `D_OPR2_RS2))))
                dbg_cntr_dep_raw <= dbg_cntr_dep_raw + 1;
            else if ((dec0_ix_rd == dec1_ix_rd) && dec0_ix_wb_en && dec1_ix_wb_en)
                dbg_cntr_dep_waw <= dbg_cntr_dep_waw + 1;
            if (dec0_is_branch && (!dec1_is_int && !dec1_is_md))
                if (dec1_is_ls)
                    dbg_cntr_str_brls <= dbg_cntr_str_brls + 1;
                else if (dec1_is_branch)
                    dbg_cntr_str_brbr <= dbg_cntr_str_brbr + 1;
                else
                    dbg_cntr_str_brother <= dbg_cntr_str_brother + 1;
        end
    end

    // Fencei handling
    reg im_invalidate_done, dm_flush_done;
    always @(posedge clk) begin
        if ((!rst) && (dec0_ix_valid) && (dec0_ix_fencei) &&
                (!ix_fencei_done)) begin
            im_invalidate_req <= 1'b1;
            dm_flush_req <= 1'b1;
            im_invalidate_done <= 1'b0;
            dm_flush_done <= 1'b0;
            if (im_invalidate_resp == 1'b1) begin
                im_invalidate_req <= 1'b0;
                im_invalidate_done <= 1'b1;
            end
            if (dm_flush_resp == 1'b1) begin
                dm_flush_req <= 1'b0;
                dm_flush_done <= 1'b1;
            end
            if (dm_flush_done && im_invalidate_done) begin
                ix_if_pc_override <= 1'b1;
                ix_if_new_pc <= dec0_ix_pc + 4;
                ix_fencei_done <= 1'b1;
            end
        end
        else begin
            ix_if_pc_override <= 1'b0;
            ix_if_new_pc <= 64'bx;
            ix_fencei_done <= 1'b0;
            im_invalidate_req <= 1'b0;
            dm_flush_req <= 1'b0;
        end
    end

    always @(posedge clk) begin
        if (ix_issue_ip0) begin
            ix_ip0_op <= dec0_ix_op;
            ix_ip0_option <= dec0_ix_option;
            ix_ip0_truncate <= dec0_ix_truncate;
            ix_ip0_br_type <= dec0_ix_br_type;
            ix_ip0_br_neg <= dec0_ix_br_neg;
            ix_ip0_br_offset <= dec0_ix_imm[20:0];
            ix_ip0_br_base <= br_base_dec0;
            ix_ip0_br_is_call <= dec0_ix_br_is_call;
            ix_ip0_br_is_ret <= dec0_ix_br_is_ret;
            ix_ip0_operand1 <= operand1_dec0_value;
            ix_ip0_operand2 <= operand2_dec0_value;
            ix_ip0_bp <= dec0_ix_bp;
            ix_ip0_bp_track <= dec0_ix_bp_track;
            ix_ip0_bt <= dec0_ix_bt;
            ix_ip0_wb_en <= dec0_ix_wb_en;
            ix_ip0_dst <= dec0_ix_rd;
            ix_ip0_pc <= dec0_ix_pc;
            ix_ip0_valid <= 1'b1;
        end
        else if (ix_ip0_ready || pipe_flush) begin
            ix_ip0_valid <= 1'b0;
        end
        if (ix_issue_ip1) begin
            ix_ip1_op <= dec1_ix_op;
            ix_ip1_option <= dec1_ix_option;
            ix_ip1_truncate <= dec1_ix_truncate;
            ix_ip1_br_type <= dec1_ix_br_type;
            ix_ip1_br_neg <= dec1_ix_br_neg;
            ix_ip1_br_offset <= dec1_ix_imm[20:0];
            ix_ip1_br_base <= br_base_dec1;
            ix_ip1_br_is_call <= dec1_ix_br_is_call;
            ix_ip1_br_is_ret <= dec1_ix_br_is_ret;
            ix_ip1_operand1 <= operand1_dec1_value;
            ix_ip1_operand2 <= operand2_dec1_value;
            ix_ip1_bp <= dec1_ix_bp;
            ix_ip1_bp_track <= dec1_ix_bp_track;
            ix_ip1_bt <= dec1_ix_bt;
            ix_ip1_wb_en <= dec1_ix_wb_en;
            ix_ip1_dst <= dec1_ix_rd;
            ix_ip1_pc <= dec1_ix_pc;
            ix_ip1_speculate <= (ix_issue_ip1_dec1 && dec0_is_branch && dec0_ix_valid);
            ix_ip1_valid <= 1'b1;
        end
        else if (ix_ip1_ready || pipe_flush) begin
            ix_ip1_valid <= 1'b0;
        end
        if (ix_issue_lsp) begin
            ix_lsp_base <= (ix_issue_lsp_dec0) ? operand1_dec0_value : operand1_dec1_value;
            ix_lsp_offset <= (ix_issue_lsp_dec0) ? dec0_ix_imm[11:0] : dec1_ix_imm[11:0];
            ix_lsp_source <= (ix_issue_lsp_dec0) ? operand2_dec0_value : operand2_dec1_value;
            ix_lsp_mem_sign <= (ix_issue_lsp_dec0) ? dec0_ix_mem_sign : dec1_ix_mem_sign;
            ix_lsp_mem_width <= (ix_issue_lsp_dec0) ? dec0_ix_mem_width : dec1_ix_mem_width;
            ix_lsp_wb_en <= (ix_issue_lsp_dec0) ? dec0_ix_wb_en : dec1_ix_wb_en;
            ix_lsp_dst <= (ix_issue_lsp_dec0) ? dec0_ix_rd : dec1_ix_rd;
            ix_lsp_pc <= (ix_issue_lsp_dec0) ? dec0_ix_pc : dec1_ix_pc;
            ix_lsp_speculate <= (ix_issue_lsp_dec1 && dec0_is_branch && dec0_ix_valid);
            ix_lsp_valid <= 1'b1;
        end
        else if (ix_lsp_ready || pipe_flush) begin
            ix_lsp_valid <= 1'b0;
        end
        if (ix_issue_md) begin
            ix_md_pc <= (ix_issue_md_dec0) ? dec0_ix_pc : dec1_ix_pc;
            ix_md_dst <= (ix_issue_md_dec0) ? dec0_ix_rd : dec1_ix_rd;
            ix_md_operand1 <= (ix_issue_md_dec0) ? operand1_dec0_value : operand1_dec1_value;
            ix_md_operand2 <= (ix_issue_md_dec0) ? operand2_dec0_value : operand2_dec1_value;
            ix_md_md_op <= (ix_issue_md_dec0) ? dec0_ix_md_op : dec1_ix_md_op;
            ix_md_muldiv <= (ix_issue_md_dec0) ? dec0_ix_muldiv : dec1_ix_muldiv;
            ix_md_speculate <= (ix_issue_md_dec1 && dec0_is_branch && dec0_ix_valid);
            ix_md_valid <= 1'b1;
        end
        else if (ix_md_ready || pipe_flush) begin
            ix_md_valid <= 1'b0;
        end
        // Trap waits for all preceeding instructions to complete and blocks all
        // proceeding instructions, so it shouldn't be affected by pipe flush
        if (ix_issue_trap) begin
            ix_trap_pc <= dec0_ix_pc;
            ix_trap_dst <= dec0_ix_rd;
            ix_trap_csr_op <= dec0_ix_csr_op;
            ix_trap_csr_id <= dec0_ix_imm[11:0];
            ix_trap_csr_opr <= operand1_dec0_value;
            ix_trap_mret <= dec0_ix_mret;
            ix_trap_int <= dec0_ix_intr;
            ix_trap_intexc <= `MCAUSE_EXCEPTION;
            ix_trap_cause <= dec0_ix_cause;
            ix_trap_valid <= 1'b1;
            trap_ongoing <= 1'b1;
        end
        // But this is affected by pipe flush. If the pipeline is being flushed,
        // Not handled exceptions are not valid
        else if (exc_pending && !pipe_flush) begin
            ix_trap_pc <= lsp_fault ? lsp_unaligned_epc : mmu_fault_epc;
            ix_trap_mret <= 1'b0;
            ix_trap_int <= 1'b1;
            ix_trap_intexc <= `MCAUSE_EXCEPTION;
            ix_trap_cause <=
                    (lsp_unaligned_load) ? (`MCAUSE_LMISALGN) :
                    (lsp_unaligned_store) ? (`MCAUSE_SMISALGN) :
                    (mmu_load_page_fault) ? (`MCAUSE_LPGFAULT) :
                    (mmu_store_page_fault) ? (`MCAUSE_SPGFAULT) : 4'bx;
            ix_trap_valid <= 1'b1;
            trap_ongoing <= 1'b1;
        end
        else if (int_pending && !pipe_flush) begin
            // Respond to interrupt
            ix_trap_pc <= dec0_ix_pc;
            //ix_trap_dst <= 5'bx;
            //ix_trap_csr_op <= 2'bx;
            //ix_trap_csr_id <= 12'bx;
            //ix_trap_csr_opr <= 64'bx;
            ix_trap_mret <= 1'b0;
            ix_trap_int <= 1'b1;
            ix_trap_intexc <= `MCAUSE_INTERRUPT;
            ix_trap_cause <=
                    trap_ix_ip[`MIE_MSI] ? `MCAUSE_MSI :
                    trap_ix_ip[`MIE_MTI] ? `MCAUSE_MTI :
                    trap_ix_ip[`MIE_MEI] ? `MCAUSE_MEI : 4'bx;
            ix_trap_valid <= 1'b1;
            trap_ongoing <= 1'b1;
        end
        else if (ix_trap_ready) begin
            if (ix_trap_valid) begin
                ix_trap_valid <= 1'b0;
            end
            else begin
                trap_ongoing <= 1'b0;
            end
        end

        if (rst) begin
            ix_ip0_valid <= 1'b0;
            ix_ip1_valid <= 1'b0;
            ix_lsp_valid <= 1'b0;
            ix_md_valid <= 1'b0;
            ix_trap_valid <= 1'b0;
            trap_ongoing <= 1'b0;
        end
    end
endmodule
